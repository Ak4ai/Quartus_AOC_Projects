library verilog;
use verilog.vl_types.all;
entity Aula2_vlg_check_tst is
    port(
        pin_name2       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Aula2_vlg_check_tst;
