library verilog;
use verilog.vl_types.all;
entity mic1_vlg_vec_tst is
end mic1_vlg_vec_tst;
