library verilog;
use verilog.vl_types.all;
entity Aula2_vlg_vec_tst is
end Aula2_vlg_vec_tst;
