library verilog;
use verilog.vl_types.all;
entity FULL_ADER_8BIT_vlg_vec_tst is
end FULL_ADER_8BIT_vlg_vec_tst;
