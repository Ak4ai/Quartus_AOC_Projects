library verilog;
use verilog.vl_types.all;
entity MIC1_DEF_vlg_vec_tst is
end MIC1_DEF_vlg_vec_tst;
